package counter_pkg;
	import uvm_pkg::*;

	`include "sequence.sv"
	`include "counter_monitor.sv"
	`include "driver.sv" 
	`include "counter_agent.sv"      
	`include "counter_scoreboard.sv"      
	`include "counter_config.sv"   
	`include "counter_env.sv"      
	`include "counter_test.sv"      
endpackage: simpleadder_pkg


