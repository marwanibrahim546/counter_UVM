class counter_configuration extends uvm_object;
	`uvm_object_utils(counter_configuration)

	function new(string name = "counter_configuration");
		super.new(name);
	endfunction: new
endclass: simpleadder_configuration 
